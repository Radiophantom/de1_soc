
module top (
  input         rst_n_i,
  input         clk_i,

  output  [7:0] led_o
);

endmodule

